[aimspice]
[description]
257
NAND Gate TR
M1 4 1 3 3 ptype l=0.25u,w=0.25u
M2 4 2 3 3 ptype l=0.25u,w=0.25u
M3 4 1 6 6 ntype l=0.25u,w=0.25u
M4 6 2 0 0 ntype l=0.25u,w=0.25u
.model ntype nmos
.model ptype pmos
VDD 3 0 DC 5V
VIN1 1 0 pulse(0 5V 0 1ns 1ns 2us 4us)
VIN2 2 0 DC 5V
[tran]
0.01
5u
X
X
0
[ana]
4 1
0
1 1
1 1 0 6
3
Time
v(4)
v(1)
[end]
