[aimspice]
[description]
146
CMOS Inverter
M1 2 1 3 3 ptype L=0.25u,W=0.25u
M2 2 1 0 0 ntype L=0.25u,W=0.25u
.model ntype nmos
.model ptype pmos
VDD 3 0 DC 5V
VIN 1 0 DC
[dc]
1
VIN
0
5
0.01
[tran]
0.01
5u
X
X
0
[ana]
1 1
0
1 1
1 1 0 5
2
vin
v(2)
[end]
